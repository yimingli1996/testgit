`timescale 1ns / 1ps

module var_clocktest(
    input[31:0] period,
    input clkin, 








