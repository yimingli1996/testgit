`timescale 1ns / 1ps

module var_clock(




